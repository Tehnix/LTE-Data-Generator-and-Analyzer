library ieee;
use ieee.std_logic_1164.all;

entity tx_contr is
port (
);
end tx_contr;

architecture behavior of tx_contr is

end behavior;